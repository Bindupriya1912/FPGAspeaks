module or(a,b,x);
  input a,b;
  output y;
  assign y=a|b;
endmodule
