module not_1(a,y);
input a;
output y;
assign y=~a;
endmodule
